module MIDI_rom(input [6:0] addr, output [22:0] period);
	always_comb begin
	case(addr)
		'd0: period = 'h5D511A;
		'd1: period = 'h58144F;
		'd2: period = 'h5322C5;
		'd3: period = 'h4E7842;
		'd4: period = 'h4A10CB;
		'd5: period = 'h45E89B;
		'd6: period = 'h41FC25;
		'd7: period = 'h3E4810;
		'd8: period = 'h3AC931;
		'd9: period = 'h377C8B;
		'd10: period = 'h345F4E;
		'd11: period = 'h316ECF;
		'd12: period = 'h2EA88D;
		'd13: period = 'h2C0A27;
		'd14: period = 'h299162;
		'd15: period = 'h273C21;
		'd16: period = 'h250865;
		'd17: period = 'h22F44D;
		'd18: period = 'h20FE12;
		'd19: period = 'h1F2408;
		'd20: period = 'h1D6498;
		'd21: period = 'h1BBE45;
		'd22: period = 'h1A2FA7;
		'd23: period = 'h18B767;
		'd24: period = 'h175446;
		'd25: period = 'h160513;
		'd26: period = 'h14C8B1;
		'd27: period = 'h139E10;
		'd28: period = 'h128432;
		'd29: period = 'h117A26;
		'd30: period = 'h107F09;
		'd31: period = 'h0F9204;
		'd32: period = 'h0EB24C;
		'd33: period = 'h0DDF22;
		'd34: period = 'h0D17D3;
		'd35: period = 'h0C5BB3;
		'd36: period = 'h0BAA23;
		'd37: period = 'h0B0289;
		'd38: period = 'h0A6458;
		'd39: period = 'h09CF08;
		'd40: period = 'h094219;
		'd41: period = 'h08BD13;
		'd42: period = 'h083F84;
		'd43: period = 'h07C902;
		'd44: period = 'h075926;
		'd45: period = 'h06EF91;
		'd46: period = 'h068BE9;
		'd47: period = 'h062DD9;
		'd48: period = 'h05D511;
		'd49: period = 'h058144;
		'd50: period = 'h05322C;
		'd51: period = 'h04E784;
		'd52: period = 'h04A10C;
		'd53: period = 'h045E89;
		'd54: period = 'h041FC2;
		'd55: period = 'h03E481;
		'd56: period = 'h03AC93;
		'd57: period = 'h0377C8;
		'd58: period = 'h0345F4;
		'd59: period = 'h0316EC;
		'd60: period = 'h02EA88;
		'd61: period = 'h02C0A2;
		'd62: period = 'h029916;
		'd63: period = 'h0273C2;
		'd64: period = 'h025086;
		'd65: period = 'h022F44;
		'd66: period = 'h020FE1;
		'd67: period = 'h01F240;
		'd68: period = 'h01D649;
		'd69: period = 'h01BBE4;
		'd70: period = 'h01A2FA;
		'd71: period = 'h018B76;
		'd72: period = 'h017544;
		'd73: period = 'h016051;
		'd74: period = 'h014C8B;
		'd75: period = 'h0139E1;
		'd76: period = 'h012843;
		'd77: period = 'h0117A2;
		'd78: period = 'h0107F0;
		'd79: period = 'h00F920;
		'd80: period = 'h00EB24;
		'd81: period = 'h00DDF2;
		'd82: period = 'h00D17D;
		'd83: period = 'h00C5BB;
		'd84: period = 'h00BAA2;
		'd85: period = 'h00B028;
		'd86: period = 'h00A645;
		'd87: period = 'h009CF0;
		'd88: period = 'h009421;
		'd89: period = 'h008BD1;
		'd90: period = 'h0083F8;
		'd91: period = 'h007C90;
		'd92: period = 'h007592;
		'd93: period = 'h006EF9;
		'd94: period = 'h0068BE;
		'd95: period = 'h0062DD;
		'd96: period = 'h005D51;
		'd97: period = 'h005814;
		'd98: period = 'h005322;
		'd99: period = 'h004E78;
		'd100: period = 'h004A10;
		'd101: period = 'h0045E8;
		'd102: period = 'h0041FC;
		'd103: period = 'h003E48;
		'd104: period = 'h003AC9;
		'd105: period = 'h00377C;
		'd106: period = 'h00345F;
		'd107: period = 'h00316E;
		'd108: period = 'h002EA8;
		'd109: period = 'h002C0A;
		'd110: period = 'h002991;
		'd111: period = 'h00273C;
		'd112: period = 'h002508;
		'd113: period = 'h0022F4;
		'd114: period = 'h0020FE;
		'd115: period = 'h001F24;
		'd116: period = 'h001D64;
		'd117: period = 'h001BBE;
		'd118: period = 'h001A2F;
		'd119: period = 'h0018B7;
		'd120: period = 'h001754;
		'd121: period = 'h001605;
		'd122: period = 'h0014C8;
		'd123: period = 'h00139E;
		'd124: period = 'h001284;
		'd125: period = 'h00117A;
		'd126: period = 'h00107F;
		'd127: period = 'h000F92;
		default: period = 'h0;
	endcase
	end
endmodule 